library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity senoidal is
    generic (
        BITS_DATO  : natural := 12;   -- Número de bits de cada dato-valor
        N_MUESTRAS : natural := 256   -- Cantidad de muestras por período de señal
    );
    port (
        clk      : in  std_logic;
        reset    : in  std_logic;
        enable   : in  std_logic;
        seno_o   : out std_logic_vector(BITS_DATO - 1 downto 0)
    );

    -- Esta función calcula la cantidad de bits necesarios 
    -- para almacenar un número entero positivo (distinto de cero)
    function log2ceil(n: positive) return natural is
        variable result: natural := 0;   -- Valor a devolver
        variable temp: positive := n;    -- Número máximo que debe almacenar
                                         -- (no puede ser cero)
      begin
        while temp > 1 loop
          result := result + 1;
          temp := temp / 2;
        end loop;
      
        if temp > 0 then
          result := result + 1;
        end if;
      
        return result;
    end function;

end entity senoidal;

architecture senoidal_arq of senoidal is
    type lut_type is array (0 to N_MUESTRAS - 1) of std_logic_vector(BITS_DATO - 1 downto 0);
    constant lut : lut_type := (
        "100000000000", "100000110010", "100001100100", "100010010110", "100011001000", "100011111010", "100100101100", "100101011110", "100110001111", "100111000000", 
        "100111110001", "101000100010", "101001010010", "101010000010", "101010110001", "101011100000", "101100001111", "101100111101", "101101101011", "101110011000", 
        "101111000101", "101111110001", "110000011100", "110001000111", "110001110001", "110010011010", "110011000011", "110011101011", "110100010010", "110100111001", 
        "110101011111", "110110000011", "110110100111", "110111001010", "110111101101", "111000001110", "111000101110", "111001001110", "111001101100", "111010001010", 
        "111010100110", "111011000001", "111011011100", "111011110101", "111100001101", "111100100100", "111100111010", "111101001111", "111101100011", "111101110110", 
        "111110000111", "111110011000", "111110100111", "111110110101", "111111000010", "111111001101", "111111011000", "111111100001", "111111101001", "111111110000", 
        "111111110101", "111111111001", "111111111101", "111111111110", "111111111111", "111111111110", "111111111101", "111111111001", "111111110101", "111111110000", 
        "111111101001", "111111100001", "111111011000", "111111001101", "111111000010", "111110110101", "111110100111", "111110011000", "111110000111", "111101110110", 
        "111101100011", "111101001111", "111100111010", "111100100100", "111100001101", "111011110101", "111011011100", "111011000001", "111010100110", "111010001010", 
        "111001101100", "111001001110", "111000101110", "111000001110", "110111101101", "110111001010", "110110100111", "110110000011", "110101011111", "110100111001", 
        "110100010010", "110011101011", "110011000011", "110010011010", "110001110001", "110001000111", "110000011100", "101111110001", "101111000101", "101110011000", 
        "101101101011", "101100111101", "101100001111", "101011100000", "101010110001", "101010000010", "101001010010", "101000100010", "100111110001", "100111000000", 
        "100110001111", "100101011110", "100100101100", "100011111010", "100011001000", "100010010110", "100001100100", "100000110010", "100000000000", "011111001101", 
        "011110011011", "011101101001", "011100110111", "011100000101", "011011010011", "011010100001", "011001110000", "011000111111", "011000001110", "010111011101", 
        "010110101101", "010101111101", "010101001110", "010100011111", "010011110000", "010011000010", "010010010100", "010001100111", "010000111010", "010000001110", 
        "001111100011", "001110111000", "001110001110", "001101100101", "001100111100", "001100010100", "001011101101", "001011000110", "001010100000", "001001111100", 
        "001001011000", "001000110101", "001000010010", "000111110001", "000111010001", "000110110001", "000110010011", "000101110101", "000101011001", "000100111110", 
        "000100100011", "000100001010", "000011110010", "000011011011", "000011000101", "000010110000", "000010011100", "000010001001", "000001111000", "000001100111", 
        "000001011000", "000001001010", "000000111101", "000000110010", "000000100111", "000000011110", "000000010110", "000000001111", "000000001010", "000000000110", 
        "000000000010", "000000000001", "000000000000", "000000000001", "000000000010", "000000000110", "000000001010", "000000001111", "000000010110", "000000011110", 
        "000000100111", "000000110010", "000000111101", "000001001010", "000001011000", "000001100111", "000001111000", "000010001001", "000010011100", "000010110000", 
        "000011000101", "000011011011", "000011110010", "000100001010", "000100100011", "000100111110", "000101011001", "000101110101", "000110010011", "000110110001", 
        "000111010001", "000111110001", "001000010010", "001000110101", "001001011000", "001001111100", "001010100000", "001011000110", "001011101101", "001100010100", 
        "001100111100", "001101100101", "001110001110", "001110111000", "001111100011", "010000001110", "010000111010", "010001100111", "010010010100", "010011000010", 
        "010011110000", "010100011111", "010101001110", "010101111101", "010110101101", "010111011101", "011000001110", "011000111111", "011001110000", "011010100001", 
        "011011010011", "011100000101", "011100110111", "011101101001", "011110011011", "011111001101"
     );

    signal lut_index : unsigned(log2ceil(N_MUESTRAS) - 1 downto 0);
    signal dato      : std_logic_vector(BITS_DATO - 1 downto 0);
    
begin
    process (clk, reset)
    begin
        if reset = '1' then
            lut_index <= (others => '0');
            dato      <= (others => '0');
        elsif rising_edge(clk) then
            if enable = '1' then
                lut_index <= lut_index + 1;
                if lut_index = N_MUESTRAS - 1 then
                    lut_index <= (others => '0');
                end if;
                dato <= lut(to_integer(lut_index));
            end if;
        end if;
    end process;

    seno_o <= dato;
end architecture senoidal_arq;
